module runway_status();
	
endmodule // runway_status