/********************************************
Testbench of air traffic control system.

Airport description:
1)Airport contains two runways perpendicular to each other
2)Runway B faces E-W direction and Runway A faces N-S

Group Number:21

Member 1:
Name:Archit Pandey
Roll:16CO153

Member 2:
Name:Mohit Bhasi
ROll:16CO126
*********************************************/

`timescale 1ns/10ps
module testbench;

/********************************************
Inputs :
1) d-signifies direction of travel bits
   00-East,10-West,01-South,11-North
2) Clock
3) Enable pin
4) A,B-they are feedback from the current circuit
   which prevents a plane from landing on an 
   already occupied runway

Ouputs :
1) signal-signifies the output generated by
   the curcuit

Other Variables:
1) a-signifies the current state of runway a
2) b-signifies the current state of runway 
3) counta-counter for runway a, counts till 15
   and clears the runway after that
4) countb-counter for runway b, counts till 15
   and clears the runway after that
********************************************/
    reg en,clk;
    reg [1:0] d;
    wire [3:0]signal;
    runway_select runway_pick(d,clk,en,signal);             //Create an object of type runway_select
    initial 
    begin        
        clk = 1'b0;
        repeat (100)
        #10 clk = ~clk;                                     //Create clock 
    end 
    initial
    begin
        $dumpfile("output.vcd");                            //Create the vcd file
        $dumpvars(0,runway_pick);                           

//Uniform direction is maintained throught the test cases, but the frequency of inputs vary and 
//hence each time assigned runway may not be in direction of travel. As each operation of landing takes 15 seconds, 
//the outputs stay for consecutive inputs. For example : if runway A and B are full and a new plane wants to land,
//the circuit will sendout the wait signal for the next 15 seconds regardless of the number of times the circuit receives an input
// until a runway becomes free

        en = 1'b1;                                          //Enable switch is turned on to make the circuit take input
        d = 2'b00;
        en = 1'b0;                                          //Disabling the switch signifies input has been succesfully given
        #10
        $monitor("Direction: %d Signal: %d", d, signal);    //Display

        #100
        en = 1'b1;                                          //Enable switch is turned on to make the circuit take input
        d = 2'b00;
        en = 1'b0;                                          //Disabling the switch signifies input has been succesfully given
        #10
        $monitor("Direction: %d Signal: %d", d, signal);    //Display

        #100
        en = 1'b1;                                          //Enable switch is turned on to make the circuit take input
        d = 2'b00;
        en = 1'b0;                                          //Disabling the switch signifies input has been succesfully given
        #10
        $monitor("Direction: %d Signal: %d", d, signal);    //Display

//At this point all the runways are full for the next 15 seconds and the frequency of input is increased
//to show that the circuit will output the wait signal for the next 15 seconds

        #20
        en = 1'b1;                                          //Enable switch is turned on to make the circuit take input
        d = 2'b00;
        en = 1'b0;                                          //Disabling the switch signifies input has been succesfully given
        #10
        $monitor("Direction: %d Signal: %d", d, signal);    //Display

        #20
        en = 1'b1;                                          //Enable switch is turned on to make the circuit take input
        d = 2'b00;
        en = 1'b0;                                          //Disabling the switch signifies input has been succesfully given
        #10                
        $monitor("Direction: %d Signal: %d", d, signal);    //Display

        #20
        en = 1'b1;                                          //Enable switch is turned on to make the circuit take input
        d = 2'b00;
        en = 1'b0;                                          //Disabling the switch signifies input has been succesfully given
        #10
        $monitor("Direction: %d Signal: %d", d, signal);    //Display
        
    end
endmodule 