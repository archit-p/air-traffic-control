/********************************************
Dataflow modelling of air traffic control system.

Airport description:
1)Airport contains two runways perpendicular to each other
2)Runway B faces E-W direction and Runway A faces N-S

Group Number:21

Member 1:
Name:Archit Pandey
Roll:16CO153

Member 2:
Name:Mohit Bhasi
ROll:16CO126
*********************************************/

module VerilogDM_126_153(d,A,B,clk,E,signal);

/********************************************
Inputs :
1) d-signifies direction of travel bits
   00-East,10-West,01-South,11-North
2) Clock
3) Enable pin
4) A,B-they are feedback from the current circuit
   which prevents a plane from landing on an 
   already occupied runway

Ouputs :
1) signal-signifies the output generated by
   the curcuit

Other Variables:
1) a-signifies the current state of runway a
2) b-signifies the current state of runway 
3) counta-counter for runway a, counts till 15
   and clears the runway after that
4) countb-counter for runway b, counts till 15
   and clears the runway after that
********************************************/
	reg a;
	reg b;
	integer counta = 0;
	integer countb = 0;
	input [1:0]d;
	input E,clk;	
	output reg [3:0]signal;
	output reg A,B;
	always@(negedge E)
	begin

		assign a=A; 											//feedback received from previous function call used
		assign b=B;												//to compute current runway status

//Below is a boolean function that generates a 4 bit output representing the runway to land on
//1010 signifies land on a, 1011 signifies land on b, 1101 signifies wait

		assign signal[3]=1;
		assign signal[2]=a&b;
		assign signal[1]=~signal[2];
		assign signal[0]=a|(~b&~d[1]);
	end
	always@(posedge clk)
	begin
		assign countb=(signal==4'b1011)?countb+1:countb+1;		//If current landing is on B, start timer  for B
		assign B=(countb>5)?1:0;								//Hold runway B full till landing takes place
		assign countb=(countb==15)?0:countb;					//Reset counter for runway b when it reaches 15

	end	
	always@(posedge clk)
	begin
		assign counta=(signal==4'b1010)?counta+1:counta+1;		//If current landing is on A, start timer  for A
		assign A=(counta<10)?1:0;								//Hold runway A full till landing takes place
		assign counta=(counta==15)?0:counta;					//Reset counter for runway b when it reaches 15

	end
endmodule
